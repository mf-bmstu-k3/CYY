---  В этом файле приводится описание центрального устройства управления ЦУУ.
-- Оно должно формировать управляющие сигналы для ОП, РП и спроектированного ранее арифметического устройства
-- Внешними сигналами для ЦУУ являются сигналы set, по которому ЦУУ, устанавливается в исходное состояние и тактовый сигнал clk
-- Для арифметического устройства оно готовит операнды А и В, задает сор и подает сигнал начала операции sno, после их подготовки
-- Из арифметического устройства оно забирает результат,
-- для умножения это 2n-разрядное произведение, для сложения -n-разрядная сумма и двухразрядный признак результата.
-- Сигналом, подтверждающим выполнение операции в арифметическом устройстве, является сигнал конца операции sko
-- Для оперативной памяти оно формирует следующие сигналы:
-- data_in_OP [7:0] - данные для записи в ОП
-- address_OP [7:0] - адрес, для обращения к ОП
-- wr_en_OP - сигнал записи в ОП, если этот сигнал не активен ОП выполняет чтение
-- Из ОП в ЦУУ поступает сигнал 
-- data_out_OP [7:0] - данные, считанные из ОП
-- Для регистровой памяти РП ЦУУ формирует следующие сигналы 
-- data_a_RP - данные для записи в РП, через порт а
-- address_a_RP [2:0] - адрес, для обращения к RП, через порт a
-- wren_a_RP - сигнал записи через порт а в РП, если этот сигнал не активен PП выполняет чтение
-- data_b_RP - данные для записи в РП, через порт b
-- address_b_RP [2:0] - адрес, для обращения к RП, через порт b
-- wren_b_RP - сигнал записи через порт b в РП, если этот сигнал не активен PП выполняет чтение
-- q_a - данные, считываемые из РП, через порт а
-- q_b - данные, считываемые из РП, через порт b

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--use IEEE.numeric_std.all; -- добавляем библиотеку
LIBRARY work;

--LIBRARY altera_mf;

--USE altera_mf.altera_mf_components.all;

ENTITY CYY_AU_OP_RP_F IS
	GENERIC (n : INTEGER := 8); -- n параметр, задает разрядность операндов
	PORT (
		clk : IN STD_LOGIC; -- тактовый сигнал
		set : IN STD_LOGIC; --  сигнал начальной установки
		f_com : BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0); -- пока задает формат команды: 2 - УП; 1 - РР; 0 - ПР
		-- Для взаимодействия с АУ
		a : BUFFER STD_LOGIC_VECTOR (n - 1 DOWNTO 0);-- первый операнд для АУ		
		b : BUFFER STD_LOGIC_VECTOR (n - 1 DOWNTO 0);-- второй операнд для АУ		

		cop : BUFFER STD_LOGIC; --  код операции 1-умножение,0 - сложение для АУ
		sno : BUFFER STD_LOGIC; -- сигнал начала операции для АУ

		rr : BUFFER STD_LOGIC_VECTOR (2 * n - 1 DOWNTO 0);-- результат из АУ
		priznak : BUFFER STD_LOGIC_VECTOR (1 DOWNTO 0); -- признак результата из АУ
		sko : BUFFER STD_LOGIC; -- сигнал конца операции из АУ
		-- Для наблюдения внутренних сигналов во время отладки проекта
		SIGNAL RA : BUFFER STD_LOGIC_VECTOR (7 DOWNTO 0);-- регистр адреса, для адресации операнда в ОП
		SIGNAL CK : BUFFER STD_LOGIC_VECTOR (7 DOWNTO 0);-- счетчик команд, для адресации текущей команды в ОП
		SIGNAL RK : BUFFER STD_LOGIC_VECTOR (7 DOWNTO 0);-- регистр команд, для хранения текущей выполняемой команды
		s_out : OUT STD_LOGIC_VECTOR(2 DOWNTO 0); -- отладочный выход для наблюдения состояний БМК
		-- Для взаимодействия с ОП		
		data_in_OP : BUFFER STD_LOGIC_VECTOR (7 DOWNTO 0); -- данные для записи в ОП
		address_OP : BUFFER STD_LOGIC_VECTOR (7 DOWNTO 0); -- адрес, для обращения к ОП
		wr_en_OP : BUFFER STD_LOGIC; -- сигнал записи в ОП, если этот сигнал не активен, ОП выполняет чтение
		data_out_OP : BUFFER STD_LOGIC_VECTOR (7 DOWNTO 0); -- данные, считанные из ОП

		-- Для взаимодействия с РП
		--		data_a_RP    : buffer STD_LOGIC_VECTOR (7 downto 0); -- данные для записи в РП, через порт а
		address_a_RP : BUFFER STD_LOGIC_VECTOR (2 DOWNTO 0); -- адрес, для обращения к RП, через порт a
		wr_en_a_RP : BUFFER STD_LOGIC; -- сигнал записи через порт а в РП, если этот сигнал не активен PП выполняет чтение
		--		data_b_RP 	 : buffer STD_LOGIC_VECTOR (7 downto 0); -- данные для записи в РП, через порт b
		address_b_RP : BUFFER STD_LOGIC_VECTOR (2 DOWNTO 0); -- адрес, для обращения к RП, через порт b
		--		wr_en_b_RP 	 : buffer std_logic;							  -- сигнал записи через порт b в РП, если этот сигнал не активен PП выполняет чтение
		q_a : BUFFER STD_LOGIC_VECTOR (7 DOWNTO 0);-- данные из РП с порта а	
		q_b : BUFFER STD_LOGIC_VECTOR (7 DOWNTO 0) -- данные из РП с порта b
	);

END ENTITY CYY_AU_OP_RP_F;

ARCHITECTURE arch OF CYY_AU_OP_RP_F IS

	-----------------------------Декларация компонента ОП на 256 байт --------------------------------------------------------------------

	COMPONENT memory
		PORT (
			address : IN STD_LOGIC_VECTOR (7 DOWNTO 0); -- адресный вход
			clock : IN STD_LOGIC; -- тактовый вход
			data : IN STD_LOGIC_VECTOR (7 DOWNTO 0); -- вход данных
			wren : IN STD_LOGIC; -- разрешение записи
			q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0) -- выход данных 
		);
	END COMPONENT;
	---------------------------------------------------------------------------------------------------------------------------------------
	-- Следующим компонентом является память регистровая RP 
	-- Декларация компонента регистровой памяти на 8 байт
	-- Содержит два порта a и b
	-- Создан в QII версии 13.1 Как его создать, есть в методичке
	COMPONENT Ram_2port_11
		PORT (
			address_a : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- адресный вход порта а
			address_b : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- адресный вход порта b
			clock : IN STD_LOGIC; -- тактовый сигнал
			data_a : IN STD_LOGIC_VECTOR(7 DOWNTO 0); -- вход данных для записи через порт а
			data_b : IN STD_LOGIC_VECTOR(7 DOWNTO 0); -- вход данных для записи через порт b
			wren_a : IN STD_LOGIC; -- разрешение записи через порт а
			wren_b : IN STD_LOGIC; -- разрешение записи через порт b
			q_a : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); -- выходная шина порта a
			q_b : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) -- выходная шина порта b
		);
	END COMPONENT;

	----------------------------------------------------------------------------------------------------------------------------------------------------
	---- Компонент Арифметическое устройство, спроектированное ранее
	-- Взят из седьмого проекта

	COMPONENT ctrl_un_BO
		GENERIC (n : INTEGER);
		PORT (
			a : IN STD_LOGIC_VECTOR(n - 1 DOWNTO 0); -- вход первого операнда
			b : IN STD_LOGIC_VECTOR(n - 1 DOWNTO 0); -- вход второго операнда
			clk : IN STD_LOGIC; -- синхросигнал
			set : IN STD_LOGIC; -- сигнал начальной установки
			cop : IN STD_LOGIC; -- код операции 
			sno : IN STD_LOGIC; -- сигнал начала операции
			rr : OUT STD_LOGIC_VECTOR(2 * n - 1 DOWNTO 0); -- результат
			priznak : OUT STD_LOGIC_VECTOR(1 DOWNTO 0); -- признак результата
			sko : OUT STD_LOGIC -- сигнал конца операции
		);
	END COMPONENT;
	------------------------------------------------------------------------------------------------------------------------------------------------
	-- Декларация сигналов, используемых в проекте 
	TYPE state_type IS (s0, s1, s2, s3, s4, s5, s6); -- определяем состояния БМК
	SIGNAL next_state, state : state_type; -- следующее состояние, текущее состояние

	SIGNAL incr_CK : STD_LOGIC := '0';-- разрешение инкремента СК
	SIGNAL summ_CK : STD_LOGIC := '0';-- вычисление адреса перехода
	SIGNAL load_RK : STD_LOGIC := '0';-- загрузка команды
	SIGNAL load_RA : STD_LOGIC := '0';-- загрузка адреса
	SIGNAL IA : STD_LOGIC_VECTOR (7 DOWNTO 0);-- исполнительный адрес операнда в ОП 
	SIGNAL incr_RA : STD_LOGIC := '0';-- разрешение инкремента РА
	-----------------------------------------------------------------------------------

BEGIN
	-- устанавливаются экземпляры компонентов OP,RP,AU
	Comp_OP : memory
	PORT MAP(address_OP, clk, data_in_OP, wr_en_OP, data_out_OP);

	----------------------------------------------------------------------------------------------------------------

	Comp_RP : Ram_2port_11 PORT MAP(
		address_a => address_a_RP, -- RK(5 downto 3), -- адрес R1
		address_b => address_b_RP, -- RK(2 downto 0), -- адрес R2
		clock => clk,
		data_a => rr(7 DOWNTO 0), -- младшую часть результата для записи суммы
		data_b => (OTHERS => '0'), -- записывать через второй порт пока не надо
		wren_a => wr_en_a_RP, -- разрешение записи в РП 
		wren_b => '0', -- через порт b запись не выполняем
		q_a => q_a, -- для наблюдения на вд
		q_b => q_b -- для наблюдения на вд
	);

	-----------------------------------------------------------------------------------------------------------------------------
	Comp_AY : ctrl_un_BO
	GENERIC MAP
		(n => 8)
	PORT MAP(a, b, clk, set, cop, sno, rr, priznak, sko);

	-------------------------------------------------------------------------------------------
	pr_CK : PROCESS (set, clk) -- этот процесс определяет поведение счетчика команд СК

	BEGIN
		IF (set = '1') THEN
			CK <= (OTHERS => '0'); --устанавливаем в начальное состояние
		ELSIF clk'event AND clk = '1' THEN
			IF (incr_CK = '1') THEN
				CK <= CK + "00000001"; -- инкремент счетчика
			ELSIF (summ_CK = '1') THEN
				CK <= CK + (RK(5) & RK(5) & RK(5 DOWNTO 0)); -- вычисление адреса перехода
			END IF;
		END IF;
	END PROCESS pr_CK;
	---------------------------------------------------------------------------------------	 
	pr_RK : PROCESS (clk) -- этот процесс определяет поведение регистра команд
	BEGIN
		IF clk'event AND clk = '1' THEN -- по положительному фронту clk
			IF load_RK = '1' THEN -- если есть разрешение на прием команды
				RK <= data_out_OP; -- выполняется прием команды с выхода ОП
			END IF;
		END IF;
	END PROCESS pr_RK;
	---------------------------------------------------------------------------------------------
	pr_RA : PROCESS (clk)-- этот процесс описывает логику работы регистра адреса RA
	BEGIN
		IF clk'event AND clk = '1' THEN -- по положительному фронту 
			IF load_RA = '1' THEN
				RA <= IA; -- если есть разрешение, то загружаем исполнительный адрес первого операнда		
			ELSIF incr_RA = '1' THEN
				RA <= RA + 1; --инкремент адреса"00000001"
			END IF;
		END IF;
	END PROCESS pr_RA;
	------------------------------------------------------------------------------------------------
	-- Ниже приводится описание устройства управления для ЦУУ.Реализованы три формата команд ПР,РР и УП
	TS : PROCESS (clk, set) -- этот процесс определяет текущее состояние МУУ
	BEGIN
		IF set = '1' THEN
			state <= s0;
		ELSIF (rising_edge(clk)) THEN -- по положительному фронту переключаются состояния
			state <= next_state;
		END IF;
	END PROCESS TS;

	NS : PROCESS (state, set, f_com, sko, priznak) -- этот процесс определяет следующее состояние МУУ, управляющие сигналы
	BEGIN
		-- 

		CASE state IS
			WHEN s0 => -- переходы из s0

				IF (set = '0') THEN
					next_state <= s1; -- если сигнал set не активен,load_RK, incr_CK 
				ELSE
					next_state <= s0; -- иначе состояние не меняется
				END IF;
			WHEN s1 =>
				IF (f_com = "00") THEN -- если формат П-Р, то
					next_state <= s2; -- переходим в s2 в случае ПР
				ELSIF (f_com = "01") THEN
					next_state <= s3; -- переходим в s3 в случае РР
				ELSIF priznak = "10" THEN
					next_state <= s6; -- переходим в s6 в случае УП и условие пер выполнено
				ELSE
					next_state <= s0; -- иначе в s0
				END IF;
			WHEN s2 =>

				next_state <= s3; -- из s2 всегда переходим в s3 load_RA,

			WHEN s3 =>
				next_state <= s4; -- из s3 всегда переходим в s4, sno=1,summ_RA

			WHEN s4 =>

				IF (sko = '1') THEN
					IF f_com = "00" THEN
						next_state <= s5; -- для формата ПР  из s4 переходим в s5, если есть sko, запись младшей части результата в ОП
					ELSE
						next_state <= s0; -- переходим в s0 для формата РР
					END IF;
				ELSE
					next_state <= s4; -- ждем завершения операции
				END IF;
			WHEN s5 =>
				next_state <= s6; -- Запись старшей части результата в ОП
			WHEN s6 =>
				next_state <= s0; -- из s6 всегда переходим в s0, это пустой такт, чтобы завершить запись в ОП и подать СК на адресный вход ОП,для выборки след ком
		END CASE;
	END PROCESS NS;
	---------------------------------------------------------------------------------------------------------
	-- ниже приводится описание управляющих сигналов для БМК

	incr_CK <= '1' WHEN (state = s0 OR (state = s1 AND f_com = "00")) ELSE -- разрешение на инкремент СК	всегда в s0  и в s1, если формат П-Р
		'0';
	summ_CK <= '1' WHEN state = s1 AND f_com = "10" AND priznak = "10" ELSE -- разрешение на приращение СК если выполняется условие перехода
		'0';
	load_RK <= '1' WHEN (state = s0) ELSE -- загрузка команды в RK всегда в s0 для любой операции
		'0';
	load_RA <= '1' WHEN (state = s2) ELSE -- загрузка ИА в RA в s2 для операции умножения
		'0';
	incr_RA <= '1' WHEN (state = s4 AND sko = '1') ELSE -- инкремент RA для записи старшей части результата в ОП, только для умножения
		'0';
	sno <= '1' WHEN (state = s3) ELSE -- когда извлекли операнды на шину А и В 
		'0';
	wr_en_OP <= '1' WHEN ((state = s4 AND sko = '1' AND f_com = "00") OR state = s5) ELSE -- запись в ОП, если П-Р 
		'0';
	data_in_OP <= rr(2 * n - 1 DOWNTO n) WHEN (state = s5) ELSE
		rr(n - 1 DOWNTO 0);

	address_OP <= CK WHEN (state = s0 OR state = s1 OR state = s6 OR f_com = "01") ELSE -- если РР, то всегда CK
		IA WHEN state = s2 ELSE
		RA;

	IA <= data_out_OP + q_a; -- вычисляем исполнительный адрес первого операнда
	wr_en_a_RP <= '1' WHEN state = s4 AND sko = '1' AND f_com = "01" ELSE -- запись в РП, если формат Р-Р
		'0';
	a <= data_out_OP WHEN f_com = "00" ELSE --на шину А- первого операнда подаем первый операнд с выхода ОП, если формат память регистр
		q_a; -- 	либо с РП с выхода данных первого порта а, если формат регистр регистр 			  
	b <= q_b; --на шину В - второго операнда подаем второй операнд, считанный через порт b РП	

	-- сигнал f_com привязываем к полю сор, задаваемому в разрядах RK[7..6]
	-- используем такое кодирование, как в восьмом проекте АУ: 00- сложение, 01-умножение
	f_com <= "00" WHEN RK(7 DOWNTO 6) = "01" ELSE -- если умн, то ПР
		"01" WHEN RK(7 DOWNTO 6) = "00" ELSE -- если сложение, то РР
		"10"; -- если переход

	cop <= RK(6); -- этот разряд определяет операцию в арифметическом устройстве
	---------------------------------------------------------------------------------------------------
	--wren_b_RP<='0'; задаем в карте портов
	address_a_RP <= RK (5 DOWNTO 3); -- поле R1  в команде
	--data_a_RP<= rr(7 downto 0); -- задаем в карте портов
	address_b_RP <= RK (2 DOWNTO 0); -- поле R2  в команде, 
	--data_b_RP<= (others=>'0'); -- задаем все нули в карте портов
	---------------------------------------------------------------------------------------------------

	-----------------------------------------------------------------------------------------------------
	--  отладочный выход для наблюдения текущего состояния
	s_out <= "000" WHEN state = s0 ELSE
		"001" WHEN state = s1 ELSE
		"010" WHEN state = s2 ELSE
		"011" WHEN state = s3 ELSE
		"100" WHEN state = s4 ELSE
		"101" WHEN state = s5 ELSE
		"110";
END arch;